enter - clockul placii
afisor - suma din contul selectat (cifra unitatilor la dreapta)
V10 - opreste 
U12,U11- combinatia care selecteaza una dintre cele 3 operatii: depunere, retragere, transfer (U12 bitul mai semnificativ)


